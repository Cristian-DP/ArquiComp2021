module ALU 
@(
    // Param
)

(
    // Port
);

// internal signal (wire/reg)

// flags

// Sensitive

enmodule
